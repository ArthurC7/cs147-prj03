// Name: logic.v
// Module: 
// Input: 
// Output: 
//
// Notes: Common definitions
// 
//
// Revision History:
//
// Version	Date		Who		email			note
//------------------------------------------------------------------------------------------
//  1.0     Sep 02, 2014	Kaushik Patra	kpatra@sjsu.edu		Initial creation
//------------------------------------------------------------------------------------------
//
// 64-bit two's complement
module TWOSCOMP64(Y,A);
//output list
output [63:0] Y;
//input list
input [63:0] A;

// TBD
wire [63:0] inv_res;
wire carryout;

INV64_1x1 inv64_inst(inv_res, A);
RC_ADD_SUB_64(Y, carryout, inv_res, 64'b1, 1'b0);

endmodule

// 64-bit inverter
module INV64_1x1(Y,A);
//output 
output [63:0] Y;
//input
input [63:0] A;

// TBD
genvar i; 

generate
for(i = 0; i < 64; i=i+1)
begin
	not not_inst(Y[i], A[i]);
end
endgenerate

endmodule


// 32-bit two's complement
module TWOSCOMP32(Y,A);
//output list
output [31:0] Y;
//input list
input [31:0] A;

// TBD
wire [31:0] inv_res32;
wire adder_co;

INV32_1x1 invert32_inst(inv_res32, A);
RC_ADD_SUB_32 add32_inst(Y, adder_co, inv_res32, 32'b1, 1'b0);

endmodule

// 32-bit registere +ve edge, Reset on RESET=0
module REG32(Q, D, LOAD, CLK, RESET);
output [31:0] Q;

input CLK, LOAD;
input [31:0] D;
input RESET;

// TBD

endmodule

// 1 bit register +ve edge, 
// Preset on nP=0, nR=1, reset on nP=1, nR=0;
// Undefined nP=0, nR=0
// normal operation nP=1, nR=1
module REG1(Q, Qbar, D, L, C, nP, nR);
input D, C, L;
input nP, nR;
output Q,Qbar;

// TBD

endmodule

// 1 bit flipflop +ve edge, 
// Preset on nP=0, nR=1, reset on nP=1, nR=0;
// Undefined nP=0, nR=0
// normal operation nP=1, nR=1
module D_FF(Q, Qbar, D, C, nP, nR);
input D, C;
input nP, nR;
output Q,Qbar;

// TBD

endmodule

// 1 bit D latch
// Preset on nP=0, nR=1, reset on nP=1, nR=0;
// Undefined nP=0, nR=0
// normal operation nP=1, nR=1
module D_LATCH(Q, Qbar, D, C, nP, nR);
input D, C;
input nP, nR;
output Q,Qbar;

// TBD

endmodule

// 1 bit SR latch
// Preset on nP=0, nR=1, reset on nP=1, nR=0;
// Undefined nP=0, nR=0
// normal operation nP=1, nR=1
module SR_LATCH(Q,Qbar, S, R, C, nP, nR);
input S, R, C;
input nP, nR;
output Q,Qbar;

// TBD

endmodule

// 5x32 Line decoder
module DECODER_5x32(D,I);
// output
output [31:0] D;
// input
input [4:0] I;

// TBD

endmodule

// 4x16 Line decoder
module DECODER_4x16(D,I);
// output
output [15:0] D;
// input
input [3:0] I;

// TBD
genvar i;
genvar j;
wire [7:0] decode3x8_res;
wire inv_i3_res;

not not_inst(inv_i3_res, I[3]);
DECODER_3x8 decode3x8_inst(decode3x8_res, I[2:0]);

generate
for(i=0; i < 8; i=i+1)
begin
	and_inst1(D[i], inv_i3_res, decode3x8_res[i]);
end
endgenerate

generate
for(j=0; j < 8; j=j+1)
begin
	and_inst1(D[j+8], I[3], decode3x8_res[j]);
end
endgenerate

endmodule

// 3x8 Line decoder
module DECODER_3x8(D,I);
// output
output [7:0] D;
// input
input [2:0] I;

//TBD
wire [3:0] line2x4_res;
wire i2_inv_res;

DECODER_2x4 decode_inst(line2x4_res, I[1:0]);
not not_inst1(i2_inv_res, I[2]);

and and_inst1(D[0], line2x4_res[0], i2_inv_res);
and and_inst2(D[1], line2x4_res[1], i2_inv_res);
and and_inst3(D[2], line2x4_res[2], i2_inv_res);
and and_inst4(D[3], line2x4_res[3], i2_inv_res);
and and_inst5(D[4], line2x4_res[0], I[2]);
and and_inst6(D[5], line2x4_res[1], I[2]);
and and_inst7(D[6], line2x4_res[2], I[2]);
and and_inst8(D[7], line2x4_res[3], I[2]);

endmodule

// 2x4 Line decoder
module DECODER_2x4(D,I);
// output
output [3:0] D;
// input
input [1:0] I;

// TBD
wire inv_res0;
wire inv_res1;

not not_inst1(inv_res0, I[0]);
not not_inst2(inv_res1, I[1]);

and and_inst1(D[0], inv_res1, inv_res0);
and and_inst2(D[1], inv_res1, I[0]);
and and_inst3(D[2], I[1], inv_res0);
and and_inst4(D[3], I[1], I[0]);

endmodule